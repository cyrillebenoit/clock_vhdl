----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Cyrille Benoit
-- 
-- Create Date:    13:53:32 02/24/2016 
-- Design Name: 
-- Module Name:    principal - Behavioral 
-- Project Name: projetS4
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
--use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity principal is
    Port ( 	clk1 	: in  STD_LOGIC;					  -- clock a�50MHz
			piezo 	: out  STD_LOGIC;					  -- buzzer
    		switch 	: in  STD_LOGIC_VECTOR (7 downto 0);  --leviers
			button 	: in  STD_LOGIC_VECTOR (3 downto 0);  -- permet l'incrementation manuelle de l'heure
			an 	 	: out STD_LOGIC_VECTOR (3 downto 0);  -- selectionne le cadran a� utiliser
			led  	: out STD_LOGIC_VECTOR (6 downto 0); -- selectionne les segments de l'afficheur
			bin 	: out STD_LOGIC_VECTOR (7 downto 0)); -- leds
end principal;

architecture Behavioral of principal is
	
	
	--Signaux du diviseur de frequence
	signal count : std_logic_vector (25 downto 0):="00000000000000000000000000";
	signal clk : std_logic :='0';	
	
	--Signaux des compteurs
	signal usec, umin, uhour: integer range 0 to 10 :=0;
	signal dsec, dmin, dhour : integer range 0 to 6 :=0;		  
	signal sec_clk : std_logic :='0';
	signal min_clk : std_logic :='0';
	signal hour_clk : std_logic :='0';
	signal Minute : std_logic :='0';
	signal Hour : std_logic :='0';
	
	--Signaux de l'affichage
	signal value : integer range 0 to 10 :=0;
	signal cadran : integer range 0 to 4 :=1;  		  -- selectionne le cadran a� utiliser (permet de changer de cadran et de savoir ou on en est)
	signal count2 : std_logic :='0';	  
	signal test_led : std_logic_vector (7 downto 0):="00000000";
	
	--CHRONOMETRE
	signal chrono_usec,chrono_umin,chrono_dsec,chrono_dmin: integer range 0 to 10 :=0;
	signal chrono_usec2,chrono_umin2,chrono_dsec2,chrono_dmin2: integer range 0 to 10 :=0;
	signal chrono_usec3,chrono_umin3,chrono_dsec3,chrono_dmin3: integer range 0 to 10 :=1;
	signal chrono_sec_clk : std_logic :='0';
	signal chrono_min_clk : std_logic :='0';
	signal countdown_sec_clk : std_logic :='0';
	signal countdown_min_clk : std_logic :='0';
	signal countdown_hour_clk : std_logic :='0';
	signal countdown_Minute : std_logic :='0';
	signal countdown_Hour : std_logic :='0';
	signal countdown_toggle_done : std_logic :='0';
	signal chrono_permut, chrono_permut_receive : std_logic:='0';
	signal buzzer_start,buzzer_toggle : std_logic :='0';
	signal buzzer_end : integer range 0 to 4 :=0;

	signal countdown_done : std_logic:='0';
	signal chrono_toggle : std_logic :='0'; -- 0 lorsque le chronom�tre est en mode set, 1 lorsqu'il est en d�compte
	
begin
	--FS1
	--Genere une clock de 1Hz (clk) et une clock d'affichage a partir d'une clock de 50MHz (clk1)
	process(clk1) 	
	begin
		if(clk1'event and clk1='1') then
			count <=count+1;
			if (count = 24999999) then 
				clk <= not clk;
				count <= "00000000000000000000000000"; 
			end if;
		end if;
	end process;
	
	--FS7 : AVSEC
	sec_clk <= count(22) when switch(0)='0' and switch(1)='0' and (button(0)='1' or button(1)='1')
	else clk;
	
	--FS2 : Compteur de secondes
	process(sec_clk)
	begin
		if(sec_clk'event and sec_clk='1') then
			--Modification des unit�s
			if(usec=9) then
				usec<=0;
				if(dsec=5) then
					Minute<='1';
					dsec<=0;
				else
					dsec<=dsec+1;
				end if;
			else
				Minute<='0';
				usec<=usec+1;
			end if;
		end if;
	end process;
	
	--FS9 : AVMIN
	min_clk <= count(22) when (switch(0)='0' and switch(1)='0' and (button(2)='1' or button(3)='1')) or (switch(0)='1' and switch(1)='0' and (button(0)='1' or button(1)='1'))
	else Minute;
	
	--FS3 : Compteur de minutes
	process(min_clk)
	begin
		if(min_clk'event and min_clk='1') then
			
			--Modification des unit�s
			if(umin=9) then
				umin<=0;
				if(dmin=5) then
					dmin<=0;
					Hour<='1';
				else
					dmin<=dmin+1;
				end if;
			else
				Hour<='0';
				umin<=umin+1;
			end if;
		end if;
	end process;
	
	--FS10 : AVHOUR
	hour_clk <= count(22) when switch(0)='1' and switch(1)='0' and (button(2)='1' or button(3)='1')
	else Hour;
	
	--FS4 : Compteur des heures
	process(hour_clk)
	begin
		if(hour_clk'event and hour_clk='1') then
			--Modification des unit�s
			if(uhour=9) then
				uhour<=0;
				dhour<=dhour+1;
			elsif(uhour=3 and dhour=2) then
				uhour<=0;
				dhour<=0;
			else
				uhour<=uhour+1;
			end if;
		end if;
	end process;
	
	--Affichage
	count2<=count(15);
	
	--Choix du cadran selon count2
	process(count2)
	begin
		if(count2'event and count2='1') then
			if(cadran=4) then
				cadran<=1;
			else
				cadran<=cadran+1;
			end if;
		end if;
	end process;
	
	--FS5 : Multiplexeur : Choix de la valeur de value � afficher en fonction des differents param�tres
	
	-- Mode MM:SS
	value <= usec when cadran=1 and switch(0)='0' and switch(1)='0' 
	else dsec when  cadran=2 and switch(0)='0' and switch(1)='0' 
	else umin when  cadran=3 and switch(0)='0' and switch(1)='0' 
	else dmin when  cadran=4 and switch(0)='0' and switch(1)='0' 

	-- Mode HH:MM
	else umin when cadran=1 and switch(0)='1' and switch(1)='0' 
	else dmin when  cadran=2 and switch(0)='1' and switch(1)='0' 
	else uhour when  cadran=3 and switch(0)='1' and switch(1)='0' 
	else dhour when  cadran=4 and switch(0)='1' and switch(1)='0' 
	
	-- Mode chrono
	else chrono_usec when cadran=1 and switch(1)='1' 
	else chrono_dsec when cadran=2 and switch(1)='1'
	else chrono_umin when cadran=3 and switch(1)='1'
	else chrono_dmin when cadran=4 and switch(1)='1';
	
	-- Convertisseur 7 segments : traduit la valeur de value en segments � afficher	
	led<="1000000"	when value=0
	else "1111001" when value=1
	else "0100100"	when value=2
	else "0110000"	when value=3
	else "0011001"	when value=4
	else "0010010"	when value=5
	else "0000010"	when value=6
	else "1111000" when value=7
	else "0000000" when value=8
	else "0010000"	when value=9
	else "0001000" when value=10	
	else "1000000";
	
	--FS6 : D�multiplexeur : Choix du cadran
	--Mode chrono set
	an <="1111" when chrono_toggle='0' and clk='0' and switch(1)='1'
	--Mode normal et chrono d�compte
	else "1110" when cadran=1
	else "1101" when cadran=2
	else "1011" when cadran=3
	else "0111" when cadran=4;
			
	--BONUS
	-- Chronom�tre
	-- Alarme
	-- Mode am/pm
	
	--FSB1 Test
	process(usec)
	begin
		-- TEST
		bin <= switch;
	end process;
	
	--Chronom�tre
	
	--FSB1
	chrono_usec <= 0 when switch(1)='1' and button(3)='1' --RESET
	else chrono_usec2 when chrono_toggle='0' --SET
	else chrono_usec3 when chrono_toggle='1'; --DECOMPTE
	
	chrono_dsec <= 0 when switch(1)='1' and button(3)='1' --RESET
	else chrono_dsec2 when chrono_toggle='0' --SET
	else chrono_dsec3 when chrono_toggle='1'; --DECOMPTE
	
	chrono_umin <= 0 when switch(1)='1' and button(3)='1' --RESET
	else chrono_umin2 when chrono_toggle='0' --SET
	else chrono_umin3 when chrono_toggle='1'; --DECOMPTE
	
	chrono_dmin <= 0 when switch(1)='1' and button(3)='1' --RESET
	else chrono_dmin2 when chrono_toggle='0' --SET
	else chrono_dmin3 when chrono_toggle='1'; --DECOMPTE
	
	
	--FSB2 : AVSEC CHRONO
	chrono_sec_clk <= count(22) when switch(1)='1' and button(0)='1' and chrono_toggle='0'
	else '0';
	
	--FSB3 : Compteur de secondes du chrono
	process(chrono_sec_clk)
	begin
		if(chrono_sec_clk'event and chrono_sec_clk='1') then
			--Modification des unit�s
			if(chrono_usec2=9) then
				chrono_usec2<=0;
				if(chrono_dsec2=5) then
					chrono_dsec2<=0;
				else
					chrono_dsec2<=chrono_dsec2+1;
				end if;
			else
				chrono_usec2<=chrono_usec2+1;
			end if;
		end if;
		if(button(3)='1') then
			chrono_usec2<=0;
			chrono_dsec2<=0;
		end if;
	end process;
	
	--FSB2 : AVMIN CHRONO
	chrono_min_clk <= count(22) when switch(1)='1' and button(1)='1' and chrono_toggle='0'
	else '0';
	
	--FSB3 : Compteur de minutes du chrono
	process(chrono_min_clk)
	begin
		if(chrono_min_clk'event and chrono_min_clk='1') then
			--Modification des unit�s
			if(chrono_umin2=9) then
				chrono_umin2<=0;
				if(chrono_dmin2=5) then
					chrono_dmin2<=0;
				else
					chrono_dmin2<=chrono_dmin2+1;
				end if;
			else
				chrono_umin2<=chrono_umin2+1;
			end if;
		end if;
		if(button(3)='1') then
			chrono_umin2<=0;
			chrono_dmin2<=0;
		end if;
	end process;
	
	--Variable d'incr�mentation des valeurs lorsque basculement en decompte
	process(chrono_toggle)
	begin
		if(chrono_toggle'event and chrono_toggle='1') then
			chrono_permut<='1';
		end if;
		if(chrono_permut_receive='1') then
			chrono_permut<='0';
		end if;
	end process;
	
	--FSB6 : Changement d'�tat du chrono
	
	process(chrono_toggle,button,switch,countdown_done)
	begin
		if(button(2)='1' and switch(1)='1') then
			chrono_toggle<='1';
		elsif((button(3)='1' and switch(1)='1') or countdown_done='1') then
			chrono_toggle<='0';
			countdown_toggle_done<='1';
			--AJOUTER PIEZO
		else
			countdown_toggle_done<='0';
		end if;
	end process;
	
	--FSB7 : AVSEC DECOMPT
	countdown_sec_clk <= clk when chrono_toggle<='1'
	else '0';
	
	
	--FSB8 : D�compteur de secondes du chrono
	process(countdown_sec_clk,chrono_permut)
	begin
		if(countdown_sec_clk'event and countdown_sec_clk='1') then
			if(chrono_usec3=0) then
				chrono_usec3<=9;
				if(chrono_dsec3=0) then
					countdown_Minute <='1';
					chrono_dsec3<=5;
				else
					chrono_dsec3<=chrono_dsec3-1;
					countdown_Minute <='0';
				end if;
			else
				countdown_Minute <='0';
				chrono_usec3<=chrono_usec3-1;
			end if;
		end if;
		if(chrono_permut='1') then
			chrono_permut_receive<='1';
			chrono_usec3<=chrono_usec2;
			chrono_dsec3<=chrono_dsec2;
		else
			chrono_permut_receive<='0';
		end if;
		if(button(3)='1') then
			chrono_usec3<=0;
			chrono_dsec3<=0;
		end if;
	end process;
	
	--FSB5 : D�compteur de minutes du chrono
	process(countdown_Minute,chrono_permut,countdown_toggle_done)
	begin
		if(countdown_Minute'event and countdown_Minute='1') then
			if(chrono_umin3=0) then
				chrono_umin3<=9;
				if(chrono_dmin3=0) then
					chrono_dmin3<=0;
					chrono_umin3<=0;
					countdown_done<='1';
				else
					chrono_dmin3<=chrono_dmin3-1;
				end if;
			else
				chrono_umin3<=chrono_umin3-1;
			end if;
		end if;
		if(chrono_permut='1') then
			chrono_permut_receive<='1';
			chrono_umin3<=chrono_umin2;
			chrono_dmin3<=chrono_dmin2;
		else
			chrono_permut_receive<='0';
		end if;
		if(countdown_toggle_done='1') then
			countdown_done<='0';
		end if;
		if(button(3)='1') then
			chrono_umin3<=0;
			chrono_dmin3<=0;
		end if;
	end process;
	
	--Activation et desactivation du buzzer
	piezo <= clk when countdown_done='1'
	else '0' when buzzer_end =0;
	
	--Compteur du buzzer
	buzzer_start <= '1' when countdown_done='1'
	else '0' when buzzer_end=0;
	
	process(clk,buzzer_start, buzzer_end)
	begin
		if(clk'event and clk='1') then
			if(buzzer_end>0) then
				buzzer_end<=buzzer_end-1;
			end if;
		end if;
		if(buzzer_start='1' and buzzer_toggle='0') then
				buzzer_toggle<='1';
				buzzer_end<=4;
		end if;
		if(buzzer_end=0) then
		 buzzer_toggle<='0';
		end if;
	end process;
	
end Behavioral;